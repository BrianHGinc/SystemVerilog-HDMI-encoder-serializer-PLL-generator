module glyphmap ( input wire [7:0] codepoint, output wire [127:0] glyph );
assign glyph = codepoint == 8'b00000000 ? 128'h00007E42424242424242427E00000000
    : codepoint == 8'b00000001 ? 128'h00007C82AA8282BA9282827C00000000
    : codepoint == 8'b00000010 ? 128'h00007CFED6FEFEC6EEFEFE7C00000000
    : codepoint == 8'b00000011 ? 128'h000000006CFEFEFEFE7C381000000000
    : codepoint == 8'b00000100 ? 128'h0000000010387CFE7C38100000000000
    : codepoint == 8'b00000101 ? 128'h00001038381054FEFE54103800000000
    : codepoint == 8'b00000110 ? 128'h00001010387CFEFE7C10103800000000
    : codepoint == 8'b00000111 ? 128'h000000000000183C3C18000000000000
    : codepoint == 8'b00001000 ? 128'hFFFFFFFFFFFFE7C3C3E7FFFFFFFFFFFF
    : codepoint == 8'b00001001 ? 128'h00000000000018242418000000000000
    : codepoint == 8'b00001010 ? 128'hFFFFFFFFFFFFE7DBDBE7FFFFFFFFFFFF
    : codepoint == 8'b00001011 ? 128'h00001E060A1238444444443800000000
    : codepoint == 8'b00001100 ? 128'h0000384444444438107C101000000000
    : codepoint == 8'b00001101 ? 128'h00003E223E202020202020C000000000
    : codepoint == 8'b00001110 ? 128'h00007E427E4242424242424480000000
    : codepoint == 8'b00001111 ? 128'h00000010925438EE3854921000000000
    : codepoint == 8'b00010000 ? 128'h00000000C0F0FCFFFCF0C00000000000
    : codepoint == 8'b00010001 ? 128'h00000000030F3FFF3F0F030000000000
    : codepoint == 8'b00010010 ? 128'h00001038541010101054381000000000
    : codepoint == 8'b00010011 ? 128'h00002424242424242400242400000000
    : codepoint == 8'b00010100 ? 128'h00007E92929292721212121200000000
    : codepoint == 8'b00010101 ? 128'h00384440304844442418044438000000
    : codepoint == 8'b00010110 ? 128'h00000000000000007E7E7E7E00000000
    : codepoint == 8'b00010111 ? 128'h00001038541010105438107C00000000
    : codepoint == 8'b00011000 ? 128'h00001038541010101010101000000000
    : codepoint == 8'b00011001 ? 128'h00001010101010101054381000000000
    : codepoint == 8'b00011010 ? 128'h00000000000804FE0408000000000000
    : codepoint == 8'b00011011 ? 128'h00000000002040FE4020000000000000
    : codepoint == 8'b00011100 ? 128'h0000000040404040407E000000000000
    : codepoint == 8'b00011101 ? 128'h00000000002442FF4224000000000000
    : codepoint == 8'b00011110 ? 128'h00000000101038387C7CFEFE00000000
    : codepoint == 8'b00011111 ? 128'h00000000FEFE7C7C3838101000000000
    : codepoint == 8'b00100000 ? 128'h00000000000000000000000000000000
    : codepoint == 8'b00100001 ? 128'h00001010101010101000101000000000
    : codepoint == 8'b00100010 ? 128'h00242424000000000000000000000000
    : codepoint == 8'b00100011 ? 128'h00002424247E24247E24242400000000
    : codepoint == 8'b00100100 ? 128'h0010107C9290907C1212927C10100000
    : codepoint == 8'b00100101 ? 128'h0000649468081010202C524C00000000
    : codepoint == 8'b00100110 ? 128'h000018242418304A4444443A00000000
    : codepoint == 8'b00100111 ? 128'h00101010000000000000000000000000
    : codepoint == 8'b00101000 ? 128'h00000810202020202020100800000000
    : codepoint == 8'b00101001 ? 128'h00002010080808080808102000000000
    : codepoint == 8'b00101010 ? 128'h000000000024187E1824000000000000
    : codepoint == 8'b00101011 ? 128'h000000000010107C1010000000000000
    : codepoint == 8'b00101100 ? 128'h00000000000000000000101020000000
    : codepoint == 8'b00101101 ? 128'h000000000000007E0000000000000000
    : codepoint == 8'b00101110 ? 128'h00000000000000000000101000000000
    : codepoint == 8'b00101111 ? 128'h00000404080810102020404000000000
    : codepoint == 8'b00110000 ? 128'h00003C4242464A526242423C00000000
    : codepoint == 8'b00110001 ? 128'h00000818280808080808083E00000000
    : codepoint == 8'b00110010 ? 128'h00003C42420204081020407E00000000
    : codepoint == 8'b00110011 ? 128'h00003C4242021C020242423C00000000
    : codepoint == 8'b00110100 ? 128'h000002060A1222427E02020200000000
    : codepoint == 8'b00110101 ? 128'h00007E4040407C020202423C00000000
    : codepoint == 8'b00110110 ? 128'h00001C2040407C424242423C00000000
    : codepoint == 8'b00110111 ? 128'h00007E02020404080810101000000000
    : codepoint == 8'b00111000 ? 128'h00003C4242423C424242423C00000000
    : codepoint == 8'b00111001 ? 128'h00003C424242423E0202043800000000
    : codepoint == 8'b00111010 ? 128'h00000000001010000000101000000000
    : codepoint == 8'b00111011 ? 128'h00000000001010000000101020000000
    : codepoint == 8'b00111100 ? 128'h00000004081020402010080400000000
    : codepoint == 8'b00111101 ? 128'h00000000007E00007E00000000000000
    : codepoint == 8'b00111110 ? 128'h00000040201008040810204000000000
    : codepoint == 8'b00111111 ? 128'h00003C42424204080800080800000000
    : codepoint == 8'b01000000 ? 128'h00007C829EA2A2A2A69A807E00000000
    : codepoint == 8'b01000001 ? 128'h00003C424242427E4242424200000000
    : codepoint == 8'b01000010 ? 128'h00007C4242427C424242427C00000000
    : codepoint == 8'b01000011 ? 128'h00003C42424040404042423C00000000
    : codepoint == 8'b01000100 ? 128'h00007844424242424242447800000000
    : codepoint == 8'b01000101 ? 128'h00007E40404078404040407E00000000
    : codepoint == 8'b01000110 ? 128'h00007E40404078404040404000000000
    : codepoint == 8'b01000111 ? 128'h00003C424240404E4242423C00000000
    : codepoint == 8'b01001000 ? 128'h0000424242427E424242424200000000
    : codepoint == 8'b01001001 ? 128'h00003810101010101010103800000000
    : codepoint == 8'b01001010 ? 128'h00000E04040404040444443800000000
    : codepoint == 8'b01001011 ? 128'h00004244485060605048444200000000
    : codepoint == 8'b01001100 ? 128'h00004040404040404040407E00000000
    : codepoint == 8'b01001101 ? 128'h000082C6AA9292828282828200000000
    : codepoint == 8'b01001110 ? 128'h000042424262524A4642424200000000
    : codepoint == 8'b01001111 ? 128'h00003C42424242424242423C00000000
    : codepoint == 8'b01010000 ? 128'h00007C424242427C4040404000000000
    : codepoint == 8'b01010001 ? 128'h00003C424242424242424A3C02000000
    : codepoint == 8'b01010010 ? 128'h00007C424242427C5048444200000000
    : codepoint == 8'b01010011 ? 128'h00003C4240403C020242423C00000000
    : codepoint == 8'b01010100 ? 128'h0000FE10101010101010101000000000
    : codepoint == 8'b01010101 ? 128'h00004242424242424242423C00000000
    : codepoint == 8'b01010110 ? 128'h00004242424242242424181800000000
    : codepoint == 8'b01010111 ? 128'h000082828282829292AAC68200000000
    : codepoint == 8'b01011000 ? 128'h00004242242418182424424200000000
    : codepoint == 8'b01011001 ? 128'h00008282444428101010101000000000
    : codepoint == 8'b01011010 ? 128'h00007E02020408102040407E00000000
    : codepoint == 8'b01011011 ? 128'h00003820202020202020203800000000
    : codepoint == 8'b01011100 ? 128'h00004040202010100808040400000000
    : codepoint == 8'b01011101 ? 128'h00003808080808080808083800000000
    : codepoint == 8'b01011110 ? 128'h00102844000000000000000000000000
    : codepoint == 8'b01011111 ? 128'h000000000000000000000000007E0000
    : codepoint == 8'b01100000 ? 128'h10080000000000000000000000000000
    : codepoint == 8'b01100001 ? 128'h00000000003C023E4242423E00000000
    : codepoint == 8'b01100010 ? 128'h00004040407C42424242427C00000000
    : codepoint == 8'b01100011 ? 128'h00000000003C42404040423C00000000
    : codepoint == 8'b01100100 ? 128'h00000202023E42424242423E00000000
    : codepoint == 8'b01100101 ? 128'h00000000003C42427E40403C00000000
    : codepoint == 8'b01100110 ? 128'h00000E10107C10101010101000000000
    : codepoint == 8'b01100111 ? 128'h00000000003E42424242423E02023C00
    : codepoint == 8'b01101000 ? 128'h00004040407C42424242424200000000
    : codepoint == 8'b01101001 ? 128'h00001010003010101010103800000000
    : codepoint == 8'b01101010 ? 128'h00000404000C04040404040444443800
    : codepoint == 8'b01101011 ? 128'h00004040404244487048444200000000
    : codepoint == 8'b01101100 ? 128'h00003010101010101010103800000000
    : codepoint == 8'b01101101 ? 128'h0000000000FC92929292929200000000
    : codepoint == 8'b01101110 ? 128'h00000000007C42424242424200000000
    : codepoint == 8'b01101111 ? 128'h00000000003C42424242423C00000000
    : codepoint == 8'b01110000 ? 128'h00000000007C42424242427C40404000
    : codepoint == 8'b01110001 ? 128'h00000000003E42424242423E02020200
    : codepoint == 8'b01110010 ? 128'h00000000005E60404040404000000000
    : codepoint == 8'b01110011 ? 128'h00000000003E40403C02027C00000000
    : codepoint == 8'b01110100 ? 128'h00001010107C10101010100E00000000
    : codepoint == 8'b01110101 ? 128'h00000000004242424242423E00000000
    : codepoint == 8'b01110110 ? 128'h00000000004242422424181800000000
    : codepoint == 8'b01110111 ? 128'h00000000008282929292927C00000000
    : codepoint == 8'b01111000 ? 128'h00000000004242241824424200000000
    : codepoint == 8'b01111001 ? 128'h00000000004242424242423E02023C00
    : codepoint == 8'b01111010 ? 128'h00000000007E04081020407E00000000
    : codepoint == 8'b01111011 ? 128'h00000C10101020101010100C00000000
    : codepoint == 8'b01111100 ? 128'h00001010101010101010101000000000
    : codepoint == 8'b01111101 ? 128'h00003008080804080808083000000000
    : codepoint == 8'b01111110 ? 128'h0062928C000000000000000000000000
    : codepoint == 8'b01111111 ? 128'h0000000010284482828282FE00000000
    : codepoint == 8'b10000000 ? 128'h00003C42424040404042423C10102000
    : codepoint == 8'b10000001 ? 128'h00002424004242424242423E00000000
    : codepoint == 8'b10000010 ? 128'h00000810003C42427E40403C00000000
    : codepoint == 8'b10000011 ? 128'h00001824003C023E4242423E00000000
    : codepoint == 8'b10000100 ? 128'h00002424003C023E4242423E00000000
    : codepoint == 8'b10000101 ? 128'h00001008003C023E4242423E00000000
    : codepoint == 8'b10000110 ? 128'h00001824183C023E4242423E00000000
    : codepoint == 8'b10000111 ? 128'h00000000003C42404040423C10102000
    : codepoint == 8'b10001000 ? 128'h00001824003C42427E40403C00000000
    : codepoint == 8'b10001001 ? 128'h00002424003C42427E40403C00000000
    : codepoint == 8'b10001010 ? 128'h00001008003C42427E40403C00000000
    : codepoint == 8'b10001011 ? 128'h00004848003010101010103800000000
    : codepoint == 8'b10001100 ? 128'h00003048003010101010103800000000
    : codepoint == 8'b10001101 ? 128'h00002010003010101010103800000000
    : codepoint == 8'b10001110 ? 128'h2424003C4242427E4242424200000000
    : codepoint == 8'b10001111 ? 128'h1824183C4242427E4242424200000000
    : codepoint == 8'b10010000 ? 128'h0810007E404040784040407E00000000
    : codepoint == 8'b10010001 ? 128'h00000000006C12729E90906C00000000
    : codepoint == 8'b10010010 ? 128'h00007E909090FC909090909E00000000
    : codepoint == 8'b10010011 ? 128'h00001824003C42424242423C00000000
    : codepoint == 8'b10010100 ? 128'h00002424003C42424242423C00000000
    : codepoint == 8'b10010101 ? 128'h00001008003C42424242423C00000000
    : codepoint == 8'b10010110 ? 128'h00001824004242424242423E00000000
    : codepoint == 8'b10010111 ? 128'h00001008004242424242423E00000000
    : codepoint == 8'b10011000 ? 128'h00002424004242424242423E02023C00
    : codepoint == 8'b10011001 ? 128'h2424003C424242424242423C00000000
    : codepoint == 8'b10011010 ? 128'h24240042424242424242423C00000000
    : codepoint == 8'b10011011 ? 128'h00000010107C92909090927C10100000
    : codepoint == 8'b10011100 ? 128'h00001824202078202020227E00000000
    : codepoint == 8'b10011101 ? 128'h000082824428107C107C101000000000
    : codepoint == 8'b10011110 ? 128'h0000F0888888F4848E84848200000000
    : codepoint == 8'b10011111 ? 128'h00000C1210107C101010101010906000
    : codepoint == 8'b10100000 ? 128'h00000810003C023E4242423E00000000
    : codepoint == 8'b10100001 ? 128'h00000810003010101010103800000000
    : codepoint == 8'b10100010 ? 128'h00000810003C42424242423C00000000
    : codepoint == 8'b10100011 ? 128'h00000810004242424242423E00000000
    : codepoint == 8'b10100100 ? 128'h0000324C007C42424242424200000000
    : codepoint == 8'b10100101 ? 128'h324C00424262524A4642424200000000
    : codepoint == 8'b10100110 ? 128'h0038043C443C007C0000000000000000
    : codepoint == 8'b10100111 ? 128'h003844444438007C0000000000000000
    : codepoint == 8'b10101000 ? 128'h00001010001010204242423C00000000
    : codepoint == 8'b10101001 ? 128'h00000000007E40404000000000000000
    : codepoint == 8'b10101010 ? 128'h00000000007E02020200000000000000
    : codepoint == 8'b10101011 ? 128'h0020602022240810204C9204081E0000
    : codepoint == 8'b10101100 ? 128'h002060202224081022468A1E02020000
    : codepoint == 8'b10101101 ? 128'h00001010001010101010101000000000
    : codepoint == 8'b10101110 ? 128'h00000000001224489048241200000000
    : codepoint == 8'b10101111 ? 128'h00000000009048241224489000000000
    : codepoint == 8'b10110000 ? 128'h88228822882288228822882288228822
    : codepoint == 8'b10110001 ? 128'hAA55AA55AA55AA55AA55AA55AA55AA55
    : codepoint == 8'b10110010 ? 128'hEEBBEEBBEEBBEEBBEEBBEEBBEEBBEEBB
    : codepoint == 8'b10110011 ? 128'h10101010101010101010101010101010
    : codepoint == 8'b10110100 ? 128'h10101010101010F01010101010101010
    : codepoint == 8'b10110101 ? 128'h101010101010F010F010101010101010
    : codepoint == 8'b10110110 ? 128'h28282828282828E82828282828282828
    : codepoint == 8'b10110111 ? 128'h00000000000000F82828282828282828
    : codepoint == 8'b10111000 ? 128'h000000000000F010F010101010101010
    : codepoint == 8'b10111001 ? 128'h282828282828E808E828282828282828
    : codepoint == 8'b10111010 ? 128'h28282828282828282828282828282828
    : codepoint == 8'b10111011 ? 128'h000000000000F808E828282828282828
    : codepoint == 8'b10111100 ? 128'h282828282828E808F800000000000000
    : codepoint == 8'b10111101 ? 128'h28282828282828F80000000000000000
    : codepoint == 8'b10111110 ? 128'h101010101010F010F000000000000000
    : codepoint == 8'b10111111 ? 128'h00000000000000F01010101010101010
    : codepoint == 8'b11000000 ? 128'h101010101010101F0000000000000000
    : codepoint == 8'b11000001 ? 128'h10101010101010FF0000000000000000
    : codepoint == 8'b11000010 ? 128'h00000000000000FF1010101010101010
    : codepoint == 8'b11000011 ? 128'h101010101010101F1010101010101010
    : codepoint == 8'b11000100 ? 128'h00000000000000FF0000000000000000
    : codepoint == 8'b11000101 ? 128'h10101010101010FF1010101010101010
    : codepoint == 8'b11000110 ? 128'h1010101010101F101F10101010101010
    : codepoint == 8'b11000111 ? 128'h282828282828282F2828282828282828
    : codepoint == 8'b11001000 ? 128'h2828282828282F203F00000000000000
    : codepoint == 8'b11001001 ? 128'h0000000000003F202F28282828282828
    : codepoint == 8'b11001010 ? 128'h282828282828EF00FF00000000000000
    : codepoint == 8'b11001011 ? 128'h000000000000FF00EF28282828282828
    : codepoint == 8'b11001100 ? 128'h2828282828282F202F28282828282828
    : codepoint == 8'b11001101 ? 128'h000000000000FF00FF00000000000000
    : codepoint == 8'b11001110 ? 128'h282828282828EF00EF28282828282828
    : codepoint == 8'b11001111 ? 128'h101010101010FF00FF00000000000000
    : codepoint == 8'b11010000 ? 128'h28282828282828FF0000000000000000
    : codepoint == 8'b11010001 ? 128'h000000000000FF00FF10101010101010
    : codepoint == 8'b11010010 ? 128'h00000000000000FF2828282828282828
    : codepoint == 8'b11010011 ? 128'h282828282828283F0000000000000000
    : codepoint == 8'b11010100 ? 128'h1010101010101F101F00000000000000
    : codepoint == 8'b11010101 ? 128'h0000000000001F101F10101010101010
    : codepoint == 8'b11010110 ? 128'h000000000000003F2828282828282828
    : codepoint == 8'b11010111 ? 128'h28282828282828FF2828282828282828
    : codepoint == 8'b11011000 ? 128'h101010101010FF10FF10101010101010
    : codepoint == 8'b11011001 ? 128'h10101010101010F00000000000000000
    : codepoint == 8'b11011010 ? 128'h000000000000001F1010101010101010
    : codepoint == 8'b11011011 ? 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF
    : codepoint == 8'b11011100 ? 128'h0000000000000000FFFFFFFFFFFFFFFF
    : codepoint == 8'b11011101 ? 128'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0
    : codepoint == 8'b11011110 ? 128'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F
    : codepoint == 8'b11011111 ? 128'hFFFFFFFFFFFFFFFF0000000000000000
    : codepoint == 8'b11100000 ? 128'h00000000003A46444444463A00000000
    : codepoint == 8'b11100001 ? 128'h0000384444487C424242427C40404000
    : codepoint == 8'b11100010 ? 128'h00007E40404040404040404000000000
    : codepoint == 8'b11100011 ? 128'h00000000007E42424242424200000000
    : codepoint == 8'b11100100 ? 128'h00007E40201008081020407E00000000
    : codepoint == 8'b11100101 ? 128'h00000000003E44444444443800000000
    : codepoint == 8'b11100110 ? 128'h00000000004242424242467A40404000
    : codepoint == 8'b11100111 ? 128'h0000000000FE10101010100C00000000
    : codepoint == 8'b11101000 ? 128'h0000107C9292929292927C1000000000
    : codepoint == 8'b11101001 ? 128'h00003C4242425A424242423C00000000
    : codepoint == 8'b11101010 ? 128'h00003C42424242424224246600000000
    : codepoint == 8'b11101011 ? 128'h00003E10083C42424242423C00000000
    : codepoint == 8'b11101100 ? 128'h00000000007C9292927C000000000000
    : codepoint == 8'b11101101 ? 128'h000002047C8A9292A27C408000000000
    : codepoint == 8'b11101110 ? 128'h000000001E20407E40201E0000000000
    : codepoint == 8'b11101111 ? 128'h000000003C4242424242424200000000
    : codepoint == 8'b11110000 ? 128'h000000007E00007E00007E0000000000
    : codepoint == 8'b11110001 ? 128'h000000000010107C1010007C00000000
    : codepoint == 8'b11110010 ? 128'h00000020100804081020007C00000000
    : codepoint == 8'b11110011 ? 128'h00000004081020100804003E00000000
    : codepoint == 8'b11110100 ? 128'h00000C12121010101010101010101010
    : codepoint == 8'b11110101 ? 128'h10101010101010101090906000000000
    : codepoint == 8'b11110110 ? 128'h000000001010007C0010100000000000
    : codepoint == 8'b11110111 ? 128'h0000000000324C00324C000000000000
    : codepoint == 8'b11111000 ? 128'h00182424180000000000000000000000
    : codepoint == 8'b11111001 ? 128'h00000000000000181800000000000000
    : codepoint == 8'b11111010 ? 128'h00000000000000101000000000000000
    : codepoint == 8'b11111011 ? 128'h00060404040444444424140C00000000
    : codepoint == 8'b11111100 ? 128'h00003824242424000000000000000000
    : codepoint == 8'b11111101 ? 128'h0018240408103C000000000000000000
    : codepoint == 8'b11111110 ? 128'h00000000003C3C3C3C3C3C0000000000
    : codepoint == 8'b11111111 ? 128'h00000000000000000000000000000000
    : 0;
endmodule
